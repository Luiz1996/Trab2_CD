CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 13 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 10 30 70 9
0 71 1366 728
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1366 728
42991634 0
0
6 Title:
5 Name:
0
0
0
49
13 Logic Switch~
5 110 148 0 1 11
0 33
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 120 629 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 CS
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 120 716 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 OE
-7 -24 7 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 110 98 0 1 11
0 34
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 222 223 0 1 11
0 8
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 110 48 0 1 11
0 35
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 137 224 0 1 11
0 32
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 120 668 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 RD
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
5 4081~
219 326 266 0 3 22
0 6 5 7
0
0 0 96 0
4 4081
-7 -24 21 -16
3 A3C
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 10 0
1 U
3549 0 0
0
0
5 4030~
219 316 356 0 3 22
0 32 8 9
0
0 0 96 0
4 4030
-7 -24 21 -16
2 A1
0 -34 14 -26
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1124742141
65 0 0 0 4 1 12 0
1 U
7931 0 0
0
0
5 4081~
219 948 565 0 3 22
0 16 15 19
0
0 0 96 270
4 4081
-7 -24 21 -16
3 A3B
-3 -34 18 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 10 0
1 U
9325 0 0
0
0
5 4081~
219 764 570 0 3 22
0 17 15 20
0
0 0 96 270
4 4081
-7 -24 21 -16
3 A3A
-3 -34 18 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 10 0
1 U
8903 0 0
0
0
5 4081~
219 551 571 0 3 22
0 18 15 21
0
0 0 96 270
4 4081
-7 -24 21 -16
4 A27D
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 8 0
1 U
3834 0 0
0
0
14 Logic Display~
6 1020 674 0 1 2
13 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 D0
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 1021 780 0 1 2
13 2
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 D2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 1020 725 0 1 2
13 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 D1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
10 Buffer 3S~
219 986 784 0 3 22
0 12 22 2
0
0 0 96 0
7 74LS126
-24 -51 25 -43
2 A2
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 3 7 0
1 U
3874 0 0
0
0
10 Buffer 3S~
219 986 729 0 3 22
0 11 22 3
0
0 0 96 0
7 74LS126
-24 -51 25 -43
2 A3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
6671 0 0
0
0
10 Buffer 3S~
219 987 679 0 3 22
0 10 22 4
0
0 0 96 0
7 74LS126
-24 -51 25 -43
2 A4
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 1755230458
65 0 0 0 4 1 7 0
1 U
3789 0 0
0
0
5 4071~
219 952 606 0 3 22
0 27 19 12
0
0 0 96 270
4 4071
-7 -24 21 -16
4 A28C
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 9 0
1 U
4871 0 0
0
0
5 4071~
219 769 607 0 3 22
0 28 20 11
0
0 0 96 270
4 4071
-7 -24 21 -16
4 A28B
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 9 0
1 U
3750 0 0
0
0
5 4071~
219 555 611 0 3 22
0 29 21 10
0
0 0 96 270
4 4071
-7 -24 21 -16
4 A28A
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 9 0
1 U
8778 0 0
0
0
5 4081~
219 410 238 0 3 22
0 7 31 25
0
0 0 96 0
4 4081
-7 -24 21 -16
4 A27C
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 8 0
1 U
538 0 0
0
0
5 4081~
219 410 535 0 3 22
0 15 31 23
0
0 0 96 0
4 4081
-7 -24 21 -16
4 A27B
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 8 0
1 U
6843 0 0
0
0
5 4081~
219 412 372 0 3 22
0 9 31 24
0
0 0 96 0
4 4081
-7 -24 21 -16
4 A27A
-7 -34 21 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 8 0
1 U
3136 0 0
0
0
5 4081~
219 328 491 0 3 22
0 8 32 15
0
0 0 96 0
4 4081
-7 -24 21 -16
2 AB
-1 -34 13 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 6 0
1 U
5950 0 0
0
0
5 4049~
219 255 235 0 2 22
0 8 6
0
0 0 96 0
4 4049
-7 -24 21 -16
3 A2C
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 3 3 0
1 U
5670 0 0
0
0
12 D Flip-Flop~
219 895 535 0 4 9
0 33 23 48 16
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A26
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6828 0 0
0
0
12 D Flip-Flop~
219 700 534 0 4 9
0 34 23 49 17
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A25
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6735 0 0
0
0
12 D Flip-Flop~
219 493 532 0 4 9
0 35 23 50 18
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A24
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8365 0 0
0
0
5 4081~
219 957 416 0 3 22
0 36 9 39
0
0 0 96 270
4 4081
-7 -24 21 -16
2 A4
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 6 0
1 U
4132 0 0
0
0
5 4081~
219 774 421 0 3 22
0 37 9 40
0
0 0 96 270
4 4081
-7 -24 21 -16
2 A5
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 2 0
1 U
4551 0 0
0
0
5 4081~
219 560 422 0 3 22
0 38 9 41
0
0 0 96 270
4 4081
-7 -24 21 -16
2 A6
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3635 0 0
0
0
5 4071~
219 961 456 0 3 22
0 42 39 27
0
0 0 96 270
4 4071
-7 -24 21 -16
2 A7
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 5 0
1 U
3973 0 0
0
0
5 4071~
219 778 464 0 3 22
0 43 40 28
0
0 0 96 270
4 4071
-7 -24 21 -16
2 A8
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 5 0
1 U
3851 0 0
0
0
5 4071~
219 587 462 0 3 22
0 44 41 29
0
0 0 96 270
4 4071
-7 -24 21 -16
2 A9
0 -34 14 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1794086229
65 0 0 0 4 1 5 0
1 U
8383 0 0
0
0
5 4081~
219 975 291 0 3 22
0 26 7 42
0
0 0 96 270
4 4081
-7 -24 21 -16
3 A10
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9334 0 0
0
0
5 4081~
219 792 291 0 3 22
0 45 7 43
0
0 0 96 270
4 4081
-7 -24 21 -16
3 A11
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
7471 0 0
0
0
5 4081~
219 578 292 0 3 22
0 46 7 44
0
0 0 96 270
4 4081
-7 -24 21 -16
3 A12
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3334 0 0
0
0
5 4073~
219 258 707 0 4 22
0 14 30 13 22
0
0 0 96 0
4 4073
-7 -24 21 -16
2 A1
0 -34 14 -26
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
3559 0 0
0
0
12 D Flip-Flop~
219 492 362 0 4 9
0 35 24 51 38
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A15
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
984 0 0
0
0
12 D Flip-Flop~
219 699 362 0 4 9
0 34 24 52 37
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A16
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7557 0 0
0
0
12 D Flip-Flop~
219 895 362 0 4 9
0 33 24 53 36
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A17
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3146 0 0
0
0
12 D Flip-Flop~
219 894 237 0 4 9
0 33 25 54 26
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A18
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5687 0 0
0
0
12 D Flip-Flop~
219 698 239 0 4 9
0 34 25 55 45
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A19
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7939 0 0
0
0
5 4049~
219 168 236 0 2 22
0 32 5
0
0 0 96 0
4 4049
-7 -24 21 -16
3 A20
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 3 0
1 U
3308 0 0
0
0
5 4049~
219 170 668 0 2 22
0 30 47
0
0 0 96 0
4 4049
-7 -24 21 -16
3 A21
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 3 0
1 U
3408 0 0
0
0
5 4081~
219 258 659 0 3 22
0 14 47 31
0
0 0 96 0
4 4081
-7 -24 21 -16
3 A22
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
9773 0 0
0
0
12 D Flip-Flop~
219 491 237 0 4 9
0 35 25 56 46
0
0 0 4192 0
3 DFF
-10 -53 11 -45
3 A23
-10 -63 11 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
691 0 0
0
0
89
1 3 2 0 0 4224 0 15 17 0 0 2
1005 784
1001 784
1 3 3 0 0 4224 0 16 18 0 0 2
1004 729
1001 729
1 3 4 0 0 8320 0 14 19 0 0 3
1004 678
1004 679
1002 679
2 0 5 0 0 4096 0 9 0 0 62 2
302 275
189 275
1 0 6 0 0 4096 0 9 0 0 61 2
302 257
276 257
2 0 7 0 0 4096 0 39 0 0 11 2
567 270
567 257
2 0 7 0 0 0 0 38 0 0 11 2
781 269
781 257
2 0 8 0 0 4096 0 10 0 0 60 4
300 365
240 365
240 366
225 366
3 0 9 0 0 4096 0 10 0 0 21 4
349 356
357 356
357 357
364 357
3 0 7 0 0 8192 0 9 0 0 11 4
347 266
357 266
357 229
381 229
0 2 7 0 0 16512 0 0 37 15 0 6
381 229
381 240
369 240
369 257
964 257
964 269
1 3 10 0 0 4224 0 19 22 0 0 3
972 679
558 679
558 641
1 3 11 0 0 4224 0 18 21 0 0 3
971 729
772 729
772 637
3 1 12 0 0 4224 0 20 17 0 0 3
955 636
955 784
971 784
0 1 7 0 0 0 0 0 23 10 0 2
374 229
386 229
1 3 13 0 0 4224 0 3 40 0 0 2
132 716
234 716
0 1 14 0 0 4096 0 0 40 18 0 3
216 623
216 698
234 698
1 1 14 0 0 4224 0 2 48 0 0 5
132 629
216 629
216 623
234 623
234 650
2 0 9 0 0 0 0 32 0 0 21 2
763 399
763 394
2 0 9 0 0 0 0 33 0 0 21 2
549 400
549 394
2 0 9 0 0 4224 0 31 0 0 54 3
946 394
364 394
364 356
2 0 15 0 0 4096 0 12 0 0 24 2
753 548
753 543
0 2 15 0 0 8192 0 0 13 24 0 3
541 543
540 543
540 549
2 0 15 0 0 4224 0 11 0 0 52 5
937 543
447 543
447 564
369 564
369 491
1 4 16 0 0 4224 0 11 28 0 0 3
955 543
955 499
919 499
1 4 17 0 0 4224 0 12 29 0 0 3
771 548
771 498
724 498
1 4 18 0 0 4224 0 13 30 0 0 3
558 549
558 496
517 496
3 0 19 0 0 4096 0 11 0 0 45 2
946 588
946 590
3 0 20 0 0 8192 0 12 0 0 47 3
762 593
763 595
763 591
3 0 21 0 0 4096 0 13 0 0 49 2
549 594
549 595
2 0 22 0 0 4096 0 18 0 0 33 2
986 740
966 740
2 0 22 0 0 8192 0 19 0 0 33 3
987 690
987 692
962 692
4 2 22 0 0 8320 0 40 17 0 0 6
279 707
279 692
966 692
966 803
986 803
986 795
2 0 23 0 0 4096 0 30 0 0 36 2
469 514
469 535
2 0 23 0 0 0 0 29 0 0 36 2
676 516
676 535
3 2 23 0 0 4224 0 24 28 0 0 3
431 535
871 535
871 517
2 0 24 0 0 4096 0 41 0 0 39 2
468 344
468 372
2 0 24 0 0 0 0 42 0 0 39 2
675 344
675 372
3 2 24 0 0 4224 0 25 43 0 0 3
433 372
871 372
871 344
2 0 25 0 0 4096 0 49 0 0 42 2
467 219
467 238
2 0 25 0 0 0 0 45 0 0 42 2
674 221
674 238
3 2 25 0 0 4224 0 23 44 0 0 3
431 238
870 238
870 219
4 1 26 0 0 8320 0 44 37 0 0 3
918 201
982 201
982 269
3 1 27 0 0 4224 0 34 20 0 0 2
964 486
964 590
0 2 19 0 0 4224 0 0 20 0 0 2
946 595
946 590
3 1 28 0 0 4224 0 35 21 0 0 2
781 494
781 591
0 2 20 0 0 4224 0 0 21 0 0 2
763 597
763 591
3 1 29 0 0 4224 0 36 22 0 0 4
590 492
590 580
567 580
567 595
0 2 21 0 0 4224 0 0 22 0 0 2
549 602
549 595
0 2 30 0 0 8320 0 0 40 74 0 3
145 668
145 707
234 707
2 0 31 0 0 4096 0 24 0 0 55 2
386 544
375 544
1 3 15 0 0 0 0 24 26 0 0 4
386 526
385 526
385 491
349 491
2 0 31 0 0 4096 0 25 0 0 55 2
388 381
375 381
0 1 9 0 0 0 0 0 25 0 0 4
359 356
373 356
373 363
388 363
3 2 31 0 0 8320 0 48 23 0 0 4
279 659
375 659
375 247
386 247
2 0 32 0 0 4096 0 26 0 0 59 2
304 500
137 500
1 0 8 0 0 4096 0 26 0 0 60 2
304 482
225 482
1 0 32 0 0 0 0 10 0 0 59 2
300 347
137 347
1 0 32 0 0 4224 0 7 0 0 0 2
137 236
137 560
0 0 8 0 0 4224 0 0 0 63 0 2
225 235
225 560
2 0 6 0 0 4224 0 27 0 0 0 2
276 235
276 561
2 0 5 0 0 4224 0 46 0 0 0 2
189 236
189 562
1 1 8 0 0 0 0 27 5 0 0 2
240 235
222 235
1 1 32 0 0 0 0 46 7 0 0 2
153 236
137 236
1 0 33 0 0 4096 0 44 0 0 67 2
870 201
846 201
1 0 33 0 0 4096 0 43 0 0 67 2
871 326
846 326
0 1 33 0 0 4096 0 0 28 86 0 3
846 160
846 499
871 499
1 0 34 0 0 4096 0 45 0 0 70 2
674 203
657 203
1 0 34 0 0 4096 0 42 0 0 70 2
675 326
657 326
0 1 34 0 0 4096 0 0 29 87 0 3
657 109
657 498
676 498
1 0 35 0 0 4096 0 41 0 0 73 2
468 326
448 326
1 0 35 0 0 0 0 49 0 0 73 2
467 201
448 201
0 1 35 0 0 4096 0 0 30 88 0 3
448 60
448 496
469 496
1 1 30 0 0 0 0 8 47 0 0 2
132 668
155 668
4 1 36 0 0 8320 0 43 31 0 0 3
919 326
964 326
964 394
4 1 37 0 0 8320 0 42 32 0 0 3
723 326
781 326
781 399
4 1 38 0 0 8320 0 41 33 0 0 3
516 326
567 326
567 400
3 2 39 0 0 4224 0 31 34 0 0 2
955 439
955 440
3 2 40 0 0 4224 0 32 35 0 0 2
772 444
772 448
3 2 41 0 0 12416 0 33 36 0 0 4
558 445
569 445
569 446
581 446
3 1 42 0 0 4224 0 37 34 0 0 2
973 314
973 440
3 1 43 0 0 4224 0 38 35 0 0 2
790 314
790 448
3 1 44 0 0 12416 0 39 36 0 0 4
576 315
576 330
599 330
599 446
1 4 45 0 0 8320 0 38 45 0 0 3
799 269
799 203
722 203
1 4 46 0 0 8320 0 39 49 0 0 3
585 270
585 201
515 201
1 0 33 0 0 4224 0 1 0 0 0 3
110 160
965 160
965 159
1 0 34 0 0 8320 0 4 0 0 0 4
110 110
110 109
963 109
963 108
1 0 35 0 0 4224 0 6 0 0 0 2
110 60
967 60
2 2 47 0 0 4224 0 47 48 0 0 2
191 668
234 668
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 78
984 200 1004 462
994 210 1008 430
78 U
N
I
D
A
D
E 
A
R
M
A
Z
E
N
A
M
E
N
T
O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
808 696 960 720
818 704 962 720
18 CHAVE DE 3 ESTADOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
108 83 260 107
118 91 262 107
18 ENTRADA DA PALAVRA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
172 163 332 187
182 171 334 187
19 ENTRADA DE ENDERE�O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
126 598 294 622
136 606 296 622
20 ENTRADAS DE CONTROLE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
439 157 556 172
453 169 564 180
16 PRIMEIRA PALAVRA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
438 282 550 297
453 294 559 305
15 SEGUNDA PALAVRA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
440 440 557 455
454 452 565 463
16 TERCEIRA PALAVRA
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
